begin zbuffer(input clk
    input[255:0] data, input[15:0] x, input[15:0] y
);

reg[255:0] buffer_info[639:0][479:0];



endmodule